module hello;
  initial begin
    $display("Hello, world!");
    $finish;
  end
endmodule
